`include "mem_common.sv"
`include "memory.sv"
`include "mem_tx.sv"
`include "mem_gen.sv"
`include "mem_intrf.sv"
`include "mem_bfm.sv"
`include "mem_monitor.sv"
`include "mem_coverage.sv"
`include "mem_agent.sv"
`include "mem_scoreboard.sv"
`include "mem_env.sv"
`include "mem_assertion.sv"
`include "mem_tb.sv"
